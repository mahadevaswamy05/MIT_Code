//interface code
//
interface fa_if();
  logic a;
  logic b;
  logic c;
  logic sum;
  logic carry;
endinterface
